library verilog;
use verilog.vl_types.all;
entity meu_fourbits_adder_tb is
end meu_fourbits_adder_tb;
